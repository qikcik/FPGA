library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Entry_VGA is
	port (
		-- core
		in_clk_50mhz			: in std_logic;
		-- simple input
		in_keys 					: in std_logic_vector(3 downto 0);
		-- simple output
		out_buzzer 				: out std_logic							:= '0';		
		out_leds 				: out std_logic_vector(3 downto 0) 	:= (others => '0');
		-- 7seg output
		out_7seg 				: out std_logic_vector(7 downto 0) 	:= (others => '0');
		out_7segDigitSelect 	: out std_logic_vector(3 downto 0)	:= (others => '0');
		-- vga output
		out_vgaHSync			: out std_logic	:= '0';
		out_vgaVSync			: out std_logic	:= '0';
		out_vgaRGB				: out std_logic_vector(2 downto 0) := (others => '0')
	);
end Entry_VGA;

architecture behaviour of Entry_VGA is

component VgaController is
	generic (
		pixelFreq				: integer := 25_000_000;

		hSync_visibleArea	: integer := 640;
		hSync_frontPorch    : integer := 16;
		hSync_syncPulse		: integer := 96;
		hSync_backPorch     : integer := 48;

		vSync_visibleArea	: integer := 480;
		vSync_frontPorch    : integer := 10;
		vSync_syncPulse		: integer := 2;
		vSync_backPorch     : integer := 33
	);
	port (
		in_clk			: in  std_logic := '0';
		
		out_vgaRGB		: out std_logic_vector(2 downto 0) := (others => '0');
		out_vgaHSync	: out std_logic := '0';
		out_vgaVSync	: out std_logic := '0';

		out_isDisplaying	: out std_logic := '0';
		out_hPos				: out integer := 0;
		out_vPos				: out integer := 0;
		in_vgaRGB			: in  std_logic_vector(2 downto 0) := (others => '0')
	);
end component;
	
	signal isDisplaying	: std_logic := '0';
	signal hPos				: integer := 0;
	signal vPos				: integer := 0;
	
	signal position		: integer := 0;
	signal rgb			   : std_logic_vector(2 downto 0) := (others => '0');
	
	signal clk_divider 	: std_logic_vector(25 downto 0) := (others => '0'); -- 50mhz/(2^26) ~= 0.75hz
	
	constant imgR : std_logic_vector( (150*150)-1 downto 0 ) :=  "101000010001000100000000000000100000000100000000000000000010100001100010000101000010100100010101001100101101101011110101010100000111010011010000010111001101001000000000000100000100000101000000100000000000001010000000011011000000001000000101000100100010100101010111010110101010101001010101011010001001100010010000000000000000000000101000100000001000100000101010000001110100001010100010100010110100010100111101111100001010101010000011010001110010100110001001001001010000100000000100000010000101000000010000000010001000011101000000000001010010000101000100001101101010101010101001101001001000011000010101110010010110000100000000000000101000001000000011000010001000010000110110000000100000101001001010011111111011010100001110101100000100101001101001000010011001010000100100000000000000000010000010100011010001000000000000010101000000010101010100101010000100001110101010000101110101010010100000100100000101001110001011001001000100000001001000000000000101000000100010010000001110000101001010100010010101111010110100100100100110010101001010101000111010100001000011011000101001101010001000000000010000000010101000100000000001000001010010010001000011010110010111100101010100100011111101010010001000001010010010000001010001000110010100100010001000000000000111000000001000000000001101001001001010010100101011101010000000101010011101001100101010100000001001000100000000011101010001000010100010101000010010000101010100000000001010010101001000100101010101111010111000100101010101000101110111101010101100000100010010000000000101010100011001010100000101010000010101001001000101101001001101000100010100101011011010000000000000010101011011011010101010100000000010100010000000000101001101001000000100100001000101000101010101010100000101000101101010100011111111011000100000000101001010010001011011010101011000010000001111000000000000010010101011010010100100001000101010111001010001010011101110110100101010110101101101000000001001010101010111101110101010101010000010100000000000000000000100101001101001010101001000101011010110001010010101101010100010111111011100100101010000010101010101010000101011011110101000000000100000000000000000000001011100010100101010101010100100111000100000100111011111010110110110101010101010100000100101010101010111011111100101110100000100001000000000000000000001000011010110101010101010110111011110101010001011010101010100101000110010101010101000001001010010010001101010111010101100000010000010000000000000000000000000101011010101001000001010101010010101010101110110110001000110101110110111000000101010010100100110110111010101010000101001001000000000000000000000010000010001010101010111101010101101001010101101101111011000101011110011010101101000001011010101010001011011101011010010101101000101000000000000000000000001000100000010000000001010101010100010100000110011110100110110111110111110100000100100100100101010110101101010101001110001010000000000000000010000000000001000100000000000000101010100100000000000111101011101011011010101010111101000010010010110010010111011110101010100101010010101000000000000000000000000100100001001010000000010010010000100000000011111110110110110111111101101010000100101010101010100011101101010111001101011010101000000000000000000000000010100100010010000001010000010100100000000101110111010111011011010110111010000010010101010101001001101111111010100101000010001000001000000000000000000100000001101010010000001001000000010101001001011010110101110110111011101010000100100111010101010110101010110111000111111000101000000100000000100000100101001000001010000010101001010101010101101010011111110110011111101101111101000100100101010101010101101111111011010011010101000000001001000000000100001010000001010100101010101110110101101111010101010101011101110101110110101000000001010101101010100010110101101101010011110011010000000000100000000011000000000000101010001011111011011110110101111010100101001010111110111111111110001010010110101101010100110101111111010001101000100000001010000000000000001000000001101011101010110111110111111111011110101000100111101111101101010000000001001011010110101010011110111010111011110101101000000010100000001010001000000000010100111111111111111101011101110110101000010101111101111111111110000100101011011011010101010111011111101000111000001000010000000000000100010000000000101111010110111011011111111111011101100101010111110111110110110001000010010110101101010100111011111101111011000010010100000100100000010000000000000000101011111111111111111111111011110101101001011011111110111111011101000010010011110101010101011111111110111010010000000000000001000000100100010010000001111101110110110101101101101111111111010101001110111111101010101000000100101101011011101001110101101011111001000000100010101000000000100000000100100000010111111111111111111111111101111010111011110111011011111111101100000001001011011100101100111111111110101100000000000000000010100101010001010111000011111011101010101101101010101111010111011101111011111110101010110010000000110111100011010011011111111011111010000000010101000000000011010000000101100001011101111111101110111111111011111101111111011110110111111111011010000100010110111101011001111101111101011001000000010001010001000000100100111111000101101011010010111111101101101110101111011111110111111101111010101000000000010101010110101011111111111111101011000001000000000001000100000000001011100101111111111111010101101111111111101011111110111101111111011110110000000010010111111011010100111111011111111000000000110010010000100000001001011111100111111010110100111110111011010101111110111111101111111011111101010100000000010101101011001011011111110111010010000000100000000010010000000000001110100101011111111111010111011111111111011111101111111111011110101101001000000000010101111001101011110111111111101010000100011000000001000000100010110111100111110110101011110101110101110111110111111111110111111111111010100000000010001010101110010111111111110101110100000001010000000101101000000000010110101010111111111010111101111111111110111111111011111110111101101101001000000000010101111011010001111110111110101010000000100100000011010000010010111111010111101010101111011111101011011011101111111111011111101111011010100000000001001010111010101111110111101101111011000000011100001111111010010000101010100101111111110101110101111111111101101111111111111111111011101101000000000000001010101011010011111101110101110001000010001101010111110101010101011111001111110101011111011111011011101111111110111110111111011111110110100000000000101010101010101111111110101111101100000000010000100101111110100100111011100111111111101101111011111111111101011111111111111011111110110101000000000000000101011010100111111111101111110000000000101101011111111111011011011111011010110110111011010111011011111111110111011110111111011111101100100000000001001010101101111011111010111110110100000000010010010110101111101101011011101111110111011101111111111110111111111111111111101011111101101110000000100000000101010101011010111111011111000000000000010000101111111110101011011111010110111111101111011101011011101111011101111111111111110111110101000000000000001011010111111111111101101111101100000000000000101111111111111011101111111111101101111011101111111111111011111111111111111101111101011010010000000001000001010101101111011110011111100001000000000010000111111011011101111110101101111011011110111011011111011110111111010110110111011111110101000100000000001011010111111111111101101111001000000000001000100111111111110111010111101111011111110111011111110111110111111111111111111111111101101100100010100000000001010101111111111110110111100011000000000010001011111111011101111111111011110101111111101110111101111111011111111111010110101111010010001000000001010010110111110111111101011111101000001000000000000010111111111111010101111101111111010101111111101111011111110111111111110111111101111010101010010000001000001011111101111110101110100011000010000010001011111111101101111111101111011111111111010111111111110111111111011011111010110111010101010001000100000010110101111111011101111111010001000000110001000010111111111110110101111011010111011011111011011101111101111011111101101111111101101000101010010010010100010101101111111110101010001011000010001000001011111111111111101111111111111101111110111111110111101111011111111111110111101011010101010101001000000010001011111111111011111110100010010001000000000010101111111111111011111101111111011111101010111101111111111011111111011101111101101001011010101001001001010010110101111101111101000101100000011010010001111111111101101110111111111110110110111111101111011111111110110101101111010110110101010101011010000100010101111111111111110001000110001001000000001010111110111111110111111111111111111111110101110111110101111111111101101101111010101001011101010100100011010100110101010101111100000011100100000010100001111111111110101011011111011011111010111111011110111111010101011111111110101111010100101011011010011010101011111111111111010001100100110010000000100101010111110111111111111011111111111111111111110111111011111111111101010111110101010010101101101101001101011010111101101111111000100100001000000010000001111111111111010110111111111111011111101011011101010110111011110111111011011101001000101010010101010111101101111111011101100110011001100001000000000101101111111111110111110111111111111101111111110111111111111110111101011111010011101010011011010110101101101010111111011111110000001001000000001010000010111101111110101111111101101111101111011010111010110101011111101111101101010100000001001010110101010111010101111111101010101010101000001010000000001001010111111111111011111111111111111111111111011110111111101101101110110110110011001000010101010110010101110101011111011011010000110100000000001010000001111011111111101110111111111011111101110111110111101011111011111011101111001000000010100101101001010110101010111110101100000101011000001010100010000010101011011111111111111101111110111111111101110101111101011101011110110110111101000000010010101101011011111111011111101010101011011100010000101010010000110101111101111111011111111111111111101111011111010111101111110110101101010100000001001010110110101101010101111011110101110101101000001101001010000001010110111110101111111111011111111101111011110101111101110101011011010101010100000100100010010110101111011111011111010101111110111100001011100000000001011011101111111111111111111111111111111110111110101011011111101101011110101001000010100101101001110101101011110111111101111111101000100100000010010001001010111111011111111111111110111110110110110111111011101101101110101010101000100100110010101101011110110111111011110111111101111000000010010010000000110101101101110111101111111111111111111111101101101110111011010101011011010010001010001101010110110111010101111110101101111111010100010000110011000010010101111110111111111111111111111111110111111110111011010101111101011101011000100101110011010010110111110110111111111110111101110000000000001010011000010101111111101111111111111111111111111111111111101110111110101010110101101010010010101100110101011110101011110111111111111111110100000000100010001001001011111101111111110111011111011011111111011110110110101010101101011010101010001010110111011010101011110101111111111111111011010001000100010011010000011111111111111111111111111111111111011101110111101101110101110010101010011001001010101010101010101111010110111111101111101011100000100000000010010101001010111111110111111111111111111111111111111101101101011110011100101010101100100101010110110101010101110111111011110111101101111000001010001010101101011111111101111111111111111011111111111111111111011011010101101011010101101010101011011011101010101110110110111111111111110011110010101000100110110101101011111111111111011101111111101111111101110101101011011010010101010010101100101010101010101001010010110111111111111110101011111001001101010011011001011011111111111011111111111111111111011111011110111101101101010101010101010101010101010101010100010101111011010111111111011111100010010110110001111101101101111111111111111111111111111111111011101001010110110110100101010101010101010101010101010010000101111010101010110111011111010000000010000011011101110101111101111111111111110111110111111101110111101101101010101010110110101010101010100011001001000101011111010101111101111111000010001000000011111111111110111111111111111110111111111111101101011010101110101010101010101010110100101010010000101000010101010111101111111111111011000000000000000011011111101011111111111111111111111111111110111011101101110101101101011011010110101110011010101011010101010110101111110111111011101110000000000001000001111111110101111111111111111111111011110111011101010110101101110101010101110111101010000101001001101000111010011110110101111111010110000000000101010011110101111111101111011011011111101110101101110111111101111010101101101110101101011110100100100110101110101111001111111111101101111100000000000010001000111111011111111011111111111111111111111110111101101110101111101110101011101011101010010010010010110110111011101011111111111111011100000000000001001101111111111011111111111111111111111101110101101111111011110101110101111101011101111110100100100101011011101111011111111111111111111000000000000000001101011111111111011111111111011111111110111111111111111110111111111101010111101011110110100011110010101010111111101011110111101111111000000001001010001111111101111111110101111111111111111111111111101111111011101111111111111111011111111111010101001010101001110111111111011111111011110000000010000001000111101111101111111111111111111110111111110111111111011111111101111101010111110111111111010111111110111010111101111111111101111111110000000101011000010111011111111011011011101111111111111111111111110111111010111111011111111111011101110111110111101010101010111111110111111111111110000000000001000101001111111111111111111111111111011111111111111101111111111111111111111111101111111111111111010111111110111001011111111111111011111100100000000100110010101111111011111111111011111111111111011011111111111010110110111111110111111011111111111111111111100010000101011011010110111111111010000000000011000100110010111011111011111111101111111111111111111111111111111011111111111011111111011111011111111110101010010000000101110111111111010100000000000000010001000111111111011111011011111111111111111110111111101110101010111110111111111111110111111111011110100000101010001011011111111111100001000100000000100100000011111011111111111111111111011111111111111011111010101010101111110111101111111111110111111111000000000001000010101111111110100001000000000000000000000000111101110101111111011011110111111111011111101111010011111111111111111111111111111111111101010010100000000100000101110101000000000000000000000000000010011111111111011111111111111110111111111101111011001001111111110111111101111111110111101111010000001001010000010110110100000000101000000000000000000000111101111111110111111111111111111111110111101111111110111111111101111111101111111111111101111000010100000100100101101010000000000000000000000000000000001110111111111111011111111111110111111101111111110111111111111111111111111101111101111111011110000100100100101010111010000000001000000000000000000010010111111111101111111111111111111111111011110111111101101110111111101111111111111111101101111111100001001001010101010111000000001000000000000000000001010111011011111110111010111011111111011101111110111111111111111111111111111111111111111111011111111000100101001010110101100000000100000000000000000100010111111111111011111111111111011010110111111111111011111111111011111101111111101111111111111011111110001001010101011111000000000000000000000000000000000011011101111111111111111111111111111111111111111111110111111111111111111111111111111101111111111111101100101101010111110000000000000000000000000010001001111111111111101111111111111111101110111111111111101111111111111111110111111101111111101111011011110001011100111110100000000000000000000000000001000101011111110111111111011111101101111111111110111111111111111111111111111110111111011111111111111111111001010110001111110000000000000000000000000010010000111111111101110111111111111111111111011111111101111101110111110111111111111111111111111111111111100000010101111011110000000000000000000000000000001001011110111110111111111111111111111111111111101111111111111111111111111111111111110111110111111111111000000001011101111000000000000000000000000001001010110111111111111111011111111111101111111111111111111111111111111011110111111111111111111111111111111000000100111111110000000000000000000000000000000100010111111111111111011101111101111111111111111111011111111011111101111111111011111111111111111111110100000001011101111000000000000000000000000010100001001011111111110111111111101111111111101101111111111111011110111111111101111111111111111111111101111010001011111111011000001000000000000000000010100000100000101010111111111111111111110111111111111111111011111111111111011111111111101111111111111111111011100101111111111000000000000000000000000100000100010000001011111111111011111111011111101111011111111111111111111111111111011110111111111110111111111100001011111111101000000000000000000000000101010010100000100000111111111111111111111111111111111111101111111111111111111111111111111111011111011110111111100101111011111000000000000000000000000110001000001000000001111111111111101111111011111111111101111111111011111111101111011111111011111111111111101100000011111111110001000000000000000000000010010100000101000000000001111111110111111111011111011111111111111111101111111111111111111111111111111111111101001001011111111000000000000000100000000001000000000000001001001001111111111111111111111111111111101101111101111011111111101111011111111111111111111110000011111011110000101000000000000000000100000000000000000000000001111111111111111111111111111111111111111111111111101111111111111111111011010111111111101011111111111000000000001000000000000000000010100000000001000001101011111011011111111101110111111111011111111111111111111011111111111111111110110111011011111111110000001001000010000000000000000000100010000000010000100101111111101111111111111111111111111111011110111111111111111011111011111111111011001011101111110000000000000000000000000000000100001000000000000000001011111111111101011111111111011111111111111111111011111111111111011111101111111111110101111101100000000010001000100000000000000001000000000000000000100011111111111111110111101111111111110111111111111110111111111111111101111011110111011001111111100100000000000000010000000000000101011000101000100000001111101111111111111111111111111101111111101111111111111110111111011111011110111110110110011111000000000000000000000000000001010100000100000000100000000111111111111111111111111111101111111111111110111111011111111111111111100111111111011011101111000000000000000000000000000000010101010101010100001000000111111101011111110101111011111111111111111111101111111111110111110111001011111111010101101110000000000000000000000000000000000000001001000010100101000111111111110111111111111111111011101111111111111111111101111111111111111110110111101111101010100000000000000000000000000000000000001100101000000000010001111111111110111110111110111111111101111111111111011111111011111111111111111110101010101110100000000000000000000000011000000001000100000010000000000010011111111111111111011111111111111111011111101111111111111111101111110111010111111111111011101000000000000000000000001010000010010001010000100001001000111111111111111111111111111011011111111111111111111101111111111111011111111101101101101111010000000000000000000000011000100000000100000100000000000000000111111111111111111110111111111111111111111111111111011111111111111111011111111111111011111000000000000000000000000000000000000000000010000000010000101111111111111111111111111111110110111111111101111111111110110111111011111011111101111111110000000000000000000000010001010000010000000001000000000000000001111111111111111111111111111111111011111111111111011111111110111110111111111111011011111000000000000000000000000000000100000000000000000000000000000101111111111011110111111111111111101111011111111111111110111111111111111110111111111111010000000000000000000000000000000000000000000000100001000000000000101101111101111111111111111111111111111111011101111111111111111111111111111111111111111000000000000000000000000001000000010000000000000000000000000010000111011111111111110111111011111111111011111111111111111101111111101111110111111111100000000000000000000000000000000000000000000000000000000000000001000011111111111101111111111111111111111111111111111111111111111011111111111111011110100000000000000000000000000000000000000010000000000000010000000000000111111110111111111101111111011111111111111111011111011110111111111101111111111111000000000000000000000000000000000000000001000000000000000000000100000011111111111111111111111111111111111111111111111111111111111111111111111111111101001000000000000000000000000000000000000000000000000000000000000001000000111111111111111111011111111111111111111111111111111111111110111111101111010000000000000000000000000000000010000000000000000000000000000000000000010000000001111111111111111111111111111111111111111111101110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111011111111111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010010111111111111111101100101111111111111111111111111110111010100000000000000000000000000000000000000000000000010000000000000000000000000000000001010101000000101110111010010010001000011111111111111111011111101000000000000000000000000000000000000000000000000010000000000000000000010000001000010000000000000000000001000000000000000000100010101111111111110110000000000000000000000000000000000000000000000000000000010100000000000000000100000000000001010000100010000100010001000000000010001000000010101111010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000010000000000000000000000000010000000100000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000010000000000000100000000000000000000000000000000010000000000000010000000000000000000000000000000000000000001000010000000000000000000000000010000000000001010000000000010100000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000010000000000000000000000000010000000000010000000000001000000000000000000000000000000000000";
	constant imgG : std_logic_vector( (150*150)-1 downto 0 ) :=  "101101010001010101010100100010100000000000000000000000000110100001100010000101001000100000010101011101101111101111110101010100000011010011110100110111101101011010010010010100100100100100000000000000000000001010000000011011000000001010000101101101101010110101110111010100100010101001010101011010011011101011010100100100100010001010101000100000000000100000101010000001110100000010101010101010110110110110111111111100001010001000000011000001111010101110101101011101010100101000000101000000000100000000010000001010000000011101000000000001010110110101010101011101101010001000101001001001001001011010010111110011010111010101000010001001101000000000000011000010001000010000110100000000101010101101011010111111111011010100000110001000000100101001111101001011011101011010110101010000101000000000000000000011010001000100000000010101000010010101110110101110101111011110101000000001010101010010100000110101000101001110101011011011010100000101001000000000000101000000000010010000001110010101101110101011010101111010110100100100100110000100000000101000111110100101000011011010101101101110101001000000010000000010101000100000001001000101010110110101101011011111011111100101010100100001010101010010001000101011010010000001110101010110110101101010101000000000000111000000001000000000001001001011011010110101101011101010000000001010010100001000101000100000001101010101000000011111010101010110101010101010010010000101000100000010101010010101001001101101011101111110111000000001000101000101100101001010101000000101010010000000100101110101011011011101010101010101010101001001010101101101001101010110110110101011011011000000000000010100010010001010101000100000001010101010000000010111011101101010100110101011010101010101010101010101010101000100101010101011111111011010100000000001000010010001010010010101011000010101001111000000100000010110101011011010110101011010101010110101010101010111101110110110101010110101001001000000001000010101000101001010100010101010001010100000000000000101000101111101101011010101001010101011010110101011010101100010101011111111011100000101010000000100010001000000100001010100101000000010100100000000000000010011011101010100101010101010100100111000101010110111011111010110110101100000000000100000000001000100010101011110100101010100000100101000000000000010000001001011110110101010101010110111001110101010101011010101010110101000110000000000101000001001010010000001000010101010101100010110100110000000000000101001010100101011010101001000001010101010010101010101110101110000000110100000000000000000100010000100100100110101010101010000101011011001000000000100000010010010010001010101010111101010101101001010101101001110011000101011110000000000101000001011010101000001010010101001000010111101101111000000000001010000101001010100000000000000001010001010100010100000110011110100110110000000000000010000100000000000101000010101101010101001111111010000000000000100010010001010001000000000000000000101000100100000000000011101011001011010000000000000001000010010010100000010101001010000000100101011111111001001000001010101000000100100000000000000000010010010000000000000011011110110110100000000000000000000100101010101010000011101100000010001111111010101000000010001001001010100010000000000000000000010000000000000000000001110101010110000000000000000000000010000101010101001000100110100000000101011110101000011100000100100000000100000000000000000000000000000000000000000000011010110101000000000000000000000000100101010001010010101000000101000111111010101000000110000010101000100101000000000000000000000000000000000000000000010111010100000000000000001000000100100101010101010001101100100000000011111101100000011001000000100100001010000000000000000000000000000000000000000000000101011000000000000000000000000001010101101010100010100000000000010011110111010010001110100100010011000000000000000000000000000000000000000000000000000101000000000000000000000010001000000110101101010000110000010100000001111011110000111010100000100100001000000000000000000000000000000000000000000000000000000000000000000000000000000001001001000010101010001000000000010011111101101100001110100100001010000000000000000000000000000000000000000000000000000000000000000000000000000010000100001011011001010101010100001000000000111010101001010101010001000100010000000000000000000000000000000000000000000000000000000000000000000000000001000000010100100101010000000001000000100011100010111100101101101000010000000000000000000000000000000000000000000000000000000000000000000000000000000101000010010011010000010101010010101000010000110000001010010101010010100100010000000000000000000000000000000000000000000000000000000000000000000000000010000000001101001011101000000000000001000001000010100010101101010000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000001011000001000100001001000101000100000101010101011100101010000000000000000000000000000000000000000000000000000000000000000000000000000010010000000110111000010010010000000100010100001000010010111001010100011010000000000000000000000000000000000000000000000000000000000000000000000000000001010000000010010101001010000101000010000010001000001010101110101001000000100000001000000000000000000000000000000000000000000000100000000000000000000000000000000010101010010001001000001001010000011000101010010001101000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000101011001010100001000000101100001000010110010110010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010001100010000001000010000001000010000001100010001010010000000000000000000000000000000000000000000000000000000001000010000010000000000000000000000000010101011000101010100010100101000001000100111000101001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100110000101010000000000100100010101010010000101000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101010001000001010100000100000010000010110101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111010000010110001000000001011000101011101001010100000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000001010001011010000001000100000000001000010101111010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100100000010100100000101001010000101010010100100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010010100000010101000001000101000010111111010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000101100010000000000001000100010000001010011010100000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000101000000010100001000000101000000010010100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000010110000000001000101001101000000000010101010010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000100000100001000001001000101000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010101000000001000101001010000000001010100100000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000010010010000100010001011100000000110001010001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100101000000000000010001101010001000010001010000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100001000000111101010010110001010000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000010000000000100101011011010101111011010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010010100000000001011001011011010001010000010000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001001000000000010110010110110101101001010000000000100000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001010111101010111010010100000010001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100010001001001010000101110101011010010001000010000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000001000100000000000000001100010111110101010010101000000000010000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000001000010000000000000001101101110110000100101100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010001000000100101000100100111010100010010000000000000100000000000000100100000100000000000000000000000000000000000000001000000000000000000000000001001000101000000000100010111001100101010010010100000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001010010101001010010101010101000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000100001101000001010110000101000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010110100000101011010010101000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000001011000001011101010101000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001010001000000000000001010100010110111010010100000000001000000010001000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100101101000011101101010101000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000100000000000000100000101000001111110010010101000000000000000101001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101010001000101111010011011000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001001011000000011011010010100100000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000101000000100010000110011010100000000000000000010001000000000001000000001000000000000000000000000000000000000000000000000000000000010000000001000000100010000100010000010111010011010000000001000000000100001000010000000100000000100000000000000000000000000000000000000000000000000000000000000000010001001001001010101000000101010101101000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010010100100010000010001010101011011010010000000010000000001000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000100000001000001001010101010100010010101000000000100000000101010010000100100000001000000000000000000000000000000000000000000000000000000000000000010010001000010000000011010101110111010101100000000000000000010000000000000000001001000010000000000000000000000000000000000000000000000000000000000000000000100010010100001100011111010101110100101000001000000010000001000100001000000000000000000000000000000000000000000000000000000000000000000000000000001000101010100000001101001011111111011011001000000000010000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000010000000010010100001110100010111110110010101000100000010000100001000100100000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000110000000000110010011001001010000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000001000011011000010101000000010101000010100010001000100000100000010000100000000000000000000000000000000000000000000000000000000000000000000000010000100000000101000000000000100000011000010000000000000010001000000010000100000000000000000000000000000000000000000000100000000000000000000010010000101000010011001000110000000000001010001010001010001001001001001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001010000010000000000101011011100000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000100001101000111000000000000111011000010010001000000001010010010100000000000000000000000000000000000000000000000000000000000000000000000010010001000000000100110110011100000000000001101100110100100001000010001001000001001000000000000001000000000000000000000000000000000000000000000000000000000010000001010010101101101000000000000101011100001010010000000010100100000000000000000000001000010000000000100000000000000000100000000001000000000000010001000000000011100101111000000001011011011101010000100100000000100010001000000000010001000010000001000100001000000010000010001010000000000000000000000000100010010110101011010000000010101011101101001010000001000000101001000100000100000000001000000000000000001000000000000001000000000010000000000000010100010000000101111011110000000101111101111100010101010000000001000101010000010001000010100010010000010000000000000010000000100010000001000000000000000000100101010101011110000000000011010111011110010101010010000000101000000010001000010000000010000000000100000010000000010000000001000000000000000000001000000001001001101100000000000101110111111010101010010101000000001110010000000010000101010000100000100000000000100000000101010100000101000000000000000000000000100110111010000000000011011101110000100001010000010001000011010100010101010001010100010000010100000000000000000000000010100000000000000000000000000000010011010000000000000001010101010010011011001010000010101110101001001010001010101010000000000000000001000000000010010000000100000000100010000010000100001110100000000100000000101101001001101001010111000001011011010101001001010010101000000000000000000000000100000001000010010010000000000000000000000001010110000001000000000000000000000000010101110000010001001011110100100111010101101010000000000000000001000001010100100101001001000000100000000000000100000101000000000000000000000000000010010101010010000000101111110110101001010100101000000000010101000000001000000010100001000101010000000000000000000010100000000000101000000000000000000000111000101001000000101111111101010101110101000010000000000000000000101001000101010100101001010000000000000100100100001010000000000000000000000000000100001110110100100000001111101010100101010101010001000000000101001000000101000000100100010101010100000100000100100010001010000000001000000000000000000010010110110111000010010101111110100001111000000000000000101000000010100000010001011011101101111111100000000000010100010101000000000000000000000000000011010111010001001000001010111011101000001101000100010000001010010000001010001001001010101101010110111000100101000000010101100000000100000000000000000101010110101110100000000011111111000000110010010001000001101001000001000000100010101101110111111011110110001001000000010110000000000000000000000000000101010011010101100101001001011111110100001010000100100000100001010001001000010101010101011001011111111111001000000000010111100000000000000000000000000010001000111101001000000101111110100001000100001010010111001010001000000010100010101101111111101111011011110001001000111010100000000000000000000000000001000101001111100010000010011111101000101001000100100001101001010101010010010100101011011110111011111111111000000010001111110000000000000000000000000010010010111111110100000101011111110010000010011010010100110100100010000001011010101110110111111111111111100000000000111010110000000000000000000000000010101001011111010100001011011111111110101000001010000010101001011010100101001010110111110111110111111111110000000001001101111000000000000000000000000001011110110111111010011101011111111011000010101001010111111010010101001001110111010110111111111111011111111000000100111111010000000000000000000000000101010101010111011010101111010101011000101010101010000000001000101011010101011010110011011010111111111111110100000001010101111000000000000000000000000010101001001011110101110111111111101101010010100000100101011010001010101111110101011101111111111111111101111000001011111111011000001000000000000000000011101010100000101010111011111111110101010010101000000001000000101101101101101101010111001111011111111111111011000100111011011000000000000000000000000110010100010010001001101111101011010101001101000100000000100101010111011111011011011010111111111010111101101100000011101111101000000000001001000000000111110110100000100000111011111111111010100101010101010000000010110101101011111011010101010111011111011110111111000101111011111000000000000000000000000110101000001000001001011111011111100101011001010100000101011010101001011111000101011111111011111111111111101000000011111110110001000000000000000000000110111110000101000000000001111110110101101010010101000001010110110010000101111011010101011111111111011101111101001001011111111000000000000000100000000011010000000000001001000001111111110100010110101000010111101000101101101010101010101101011111101111111111010110000011111011100000101001000000000000000100001000010010000000000001111110110101010101010100000101111110110010101010101101110111101111111011010111111011100011011111111000000000001000100000000001010010100000000001000001101011101001001011100000110111011101011101010111010101011001111111110111110110110110000011111111110000001001000010000000000000001010101010000000010000100000111101101010101010111111101111010101001010110111011110101011111010111111111010000001101111110000000000000000000000000000100110101010000000000000001011101010011000010101101101011101110101101101011001101011111110010111101111010110000000111101100000000010001000100000000000010101101010100010000000000010111111100101010111101111101111010010110111101110111101011011111101101011110101000000101111100100000000000000010000000001010111011010101000100000000111101010011010101010101010101000101110101010110101010110111111011011011110111110000000011111000000000000000000000000000001011101010101010100100000000111111111001111111010110101000101001010101110110111010101011111011111100111011011000000001111000000000000000000000000000001011101111111010101001000000111110101010111110000001000100010101010110110101010110110110111110101000011110110000000000110000000000000000000000000000000000100101011010110100101000011111101010111111111100100010001001010111111101110110101010110111111111110110101000000000000000000000000000000000000000000101001011110111010010000010001111111111110111110111010010010110101010101011011011010101011111110110101010110000000000000000000000000000000000000011100001001010101001010000000000010011111111111111111011101011010110101011111101111011011010101001111110111010010100000000000000000000000000000000000001010100010010101011010100001001000111111111111111111110111011010010111011101101110110000010110110111011010101000000000000000000000000000000000000000011100101010100101000110100000000000000111111111111110111010101110111011101111111111011101000101010101101010001010000000000000010000000000000000000000000010100000001000101010000000010000001111111111111011111111111011010101111110110101110110111010100011010001010001010000000000000000000000000000000000010001010001010100000001000000000000000001111111111111011010111111011101111011111101011010001101010000010100010100000000000000000000000000000000000000000001010100000000000000000000000000000101111111111011110111111111110111101111011111111111111010101101010101101010010000000000000000000000000000000000000000000000000000000000100001000000000000101101101101110110111111111011111111111111011101011111100100101010110101010010010000010000000000000000000000000001000000010000000000000000000000000010000101011010111111110111111011111111111011111111110101011101101010100100000000000010000000000000000000000000000000010000000000000000000000000000000001000011011111111101111111111111111111111111111111111111110101011010110101010100000000000000000000000000000000000000000000000010000000000000010000000000000111110110111111111101111111011111111111111111011111011110110111010100101010001010000000000000000000000000000010000000010001000000000000000000000100000011111111111111111111111111111111111111111111111011110110111011110110110101001000001000000000000000000000000000000000000000000000000000000000000001000000111110111111111111011111111111111111111111111111111111111110011101101101000000000000000000000000000000000010100000000000100000000000000000000000010000000001111111111111111111111111111111111111111010101010111111101101101110100000000000000000000000000000000000001000000000000000000000001000000101000000000001111111111111111111111111111111111111011111111111111101011111110000000000000000000000000000000000000000000000000000000000000000000000000000100100000000010010011111111111111101100001111111111111111111101111010111000000000000000000000000000000000000000000000000001010000000000000001000000010000000001000100000000001101111000000000000000011111111111111111011111100000000000000000000000000000000000000000000010000010101000000000000000010100001010010000000000000000000000000000000000000000000010101111111111111010000000000000000000000000000000000000000000000000010101010100000000000001010101000000000001010000100010000100000001000000000000000000000010001101000000000000000000000000000000000000000000000000000000000001010100000000000000001001010100001000010000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000100100000000000000001101010000000000010000000000000100000000000000000000000000000000010000000000000010000000000000000000000000000000000000000001000010100101000000000000000001010100000000001010000000000010100000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000010000000000000001001010101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001010010000000000000000100010100000000000000000000000010000000000000000000000000010000000000010000000000001000000000000000000000000000000000000";
	constant imgB : std_logic_vector( (150*150)-1 downto 0 ) :=  "101101010000000000000000000000000000000000000000000000000110100001100010000101011010100100010101011101101111101111110001000100000011010010000000000000101101011010000000000000000000000000000000000000000000001010000000011011000000001011000101101101101010110101110111010100100010101001010000000000000000101011010100100000000000000000000000000000000000100000100010000001110100001010101010101010110111110110111111111100000000001000000011010000001000000000101101011101010100000000000000000000000100000000010000001010000000011101000000100001010110110101010101011101101000001000100001001001001001000000000000110011010111010101000000000000000000000000000011000010000000010000110110000000101110101101011010111111111010010000000100001000000100101000010000000000011101011010110101010000100000000000000000000011010001000100000000010101000010010101110111101110101111011110001000000000010001010010100000010000000000001110101011011011010100000000000000000000000101000000000010010000001110010101101110101011010101111010110100100000000010000100000000101000000000000000000011011010101101101110101001000000010000000010101000100000001001000101010110110101111011011111011111100100000000000001010101010010001000100000000000000001110101010110110101101010101000000000000111000000001000000000001101001011011010110101101011101010000000000000010000001000101000100000000000000000000000011111010101010110101010101010010010000101010100000010101010010101001001101101011101111110111000000000000100000000100001001010101100000000000000000000000101110101011011011101010101010101010101001001010101101101001101010111110110101011011011000000000000000000010000001010100000100000000000000000000000000011011101101010100110101011010101010101010101010101010101000101101010101011111111011010100000000000000000010001010010010101011000010000000100000000100000000110101011011010110101011010101010111101010101010111101110110110101010110101101000000000001000000100000000001010000010101010000000000000000000000000000101111101101011010101001010101011010110101011010101101010101011111111011100000100010000000000000001000000000001010100101000000000000000000000000000000010001001010100101010101010100100111000101010110111011111010110110111101000000000100000000000000000010000001110100101010100000000000000000000000000000001001001110110101010101010110111011110101010101011010101010110101000110000000000000000000000000000000001000000101010101100000100000000000000000000000000000000001011010101001000001010101010010101010101110111110001000110100000000000000000000000000000000100010101010001010000000000000001000000000000000000000000000001010101010111101010101101001010101101101111011000101011110000000000000000000000000001000000000010001001000000101000000000000000000000000000000000010100000000000000001010001010100010100000110011110100110110100000000000010000000000000000001000010001100010101000101010000000000000000000000000000000001000000000000000000101010100100000000000011101011101011010010000000000000000000000000000000000001001010000000100000001000000000000000000000000000000000100000000000000000010010010000100000000011011110110110100000000000000000000000000010100010000001001100000010001010100000000000000000000000000000000000000000000000000001010000010000000000000101110111010111010000000000000000000000000000010101000000000110100000000100011000001000000100000000000000000100000000000000000000000001000000000100000001011010110101000000000000000000000000000001000000010000100000000101000111010000000000000000000000000000000101000000000000000000000000000000000001000000010111110100000000000000001000000000000100010101010000100100100001000011111000000000000000000000000000001010000000000000000000000000000000000000000000010101011000000000000000000000000000000001000000000000000000000000010011100000000000000100000000000001000000000000000000000000100000000100000000000000000101001000000000000100000010000000000010101101000000100000010100000001110001000000000000000000000100000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000010001000001000000000010011101000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000100000000010000000000010001001000100000000001000000000110000000000000000000000000100010000000000000000000000000000001000000000000000000100000001000000000000000001000000000100100101010000000001000000100011100000000000000000000000000000000000000000000000000000100000000001000000000001000000000000001000000000000101000000000001010000010001010000101000010010100000000000000000000000000100010000000000100000100000000000000000000010010000000000000000000000000000000010000000000000001011100000000000000001000001000010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001000100001001000101100100000000010000001000000000000000000000000000000000000000000000000000000000000001000100000000000000000010010000000010010000010010000000000100010100011000000000010000000000011010000000100000000000000000000000000000000000000000000000000000000000000000000001010000000000010001001010000101000010000010011000000010101000000000000000100000001000000000000000000000100000000000100000000000100000000000000100000000000000000000000010010001001000001001011000011000100000000000000000100000000000000000000000000000000000000000001000000000000000000000000010000000100010000000000000001001001010000001000000101100011000000110000000000000000000000000001000001000000010000000000000000000000000100000000000000000000000000000100000000000000100010000000000010000001010011000001000000000000000000000000000000000000000000000000000000000000000000000001000010000010000000000000000000000000010000010000101010100010100101000011000000111000000000000000000000000000100000000000000000000000000000100010000000000000100000001000000000000000000000000000000100000100010000000000100101010000010000000000000000000000000000000000000000000000000000100000000000000010100000000000000000000000000000000000000000010001000001000100010100000111000000010100000010000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000101010000000110001000000001011000100000000000010100000010000000000000000000000000000000000000000000000000000100100000010000000000100000000000000001000000001010000001000100000100011000000000010000000000000000000000000000001000000000000000000000001000000000100000000001000000010000000000000000000000000000100000010100100000101001111000100000000000100100100000000010001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010100000010101000001000111000010010010000000000000000010000000000000000000000000000010000000001000000000000000000000001000000000000000000000000000001000010000000000101000110110100000000000010100000100000000000000000000000010000000000000000000000010000000001000000000000000000000000000000000000100000001000000010100001000001111000000000000000000000000000000000000000000000000000000000000000000000000001000000010000010000000000000000000000000000000000010010000000001000101001101100000000000001010010000000000000100001000000000010000000000000010000000000000000000010000000000000000000000000000000000000000000100001000001001001111000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000001000100000000000000000000001000010001000000001000101001110000000000000100110000000000000000000000000000000000010000000000000000000000100000000000100000000000000000000000000000000000000000010010000110010101111100000000100001010001000000000000000000000000000000000000100000000000010000001001000000000000000000000000000000000000000000001000000001000010001101110000000000001011010000100001000000000100000000010000000000001000000000000000000000000000000000000010000000000000000000000000001000000000100001000101111100000000100011010000001000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000100101011111010000000001011010001000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010010100000000011011000000000010001010000010000100000000100000000000000100000000000000000000000000100100100010000000000000000000000000000000000001001000100001010110111110100000000001111010000000100001000000010000001000000000000000000000000100010000000000000000000000000000000000000000000000000000000000010000000001011111100000000010011100000010001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010001001001010001111110100000000011001010010000000000000000000100001000000000000000000010000000000000000000001000000000000000000000000000000001000000000000000000001100111111110000000010111100000000010000000000000000000000100000010000000000000000000000000001000000000010000000000000000000000000001000010000000001000001111101100100000110101100000010000001000000000000000000000000000010000000000000000000001000000001000000000000000000000000001000000000001001000100101001110100110010000010111001000000100100000000000000100100000100000000000000000000010000000000000000001000000000000000000000000001001000101000000000100111111001000000000111011100000100000010000000000000000000000000000000000000000000000010000000001000000001000000000000000000000000000000001010001001010011111001000000000010111010000000100000000100100000000010000000000000000000000000000000000010000000000000000000000000000000000000000100010100000000101011101000000000000010111010000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000011110100000101000011011101000000000101000000001000000000001000000000100000100000000000100000000010000000000000000000000000000000000000001000000100000101011000000000000111111010000000000000001000000000100000000001000000000000000000000000000100000000001000000000000000000000000000001010001000000000000011010000010110010010011100000000001000000010001000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100101101000001001100111111101000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000100000000000000100010100000001111010011011101000010000000000101001000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000101010001000001011000111111101000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001001010000000001001010111100100000000000000010000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000101000000000000000000111111110000000100000000010001000000000001000000001000000000000000000000000001000000000000000000000000000000010000000001000010100010100100000000000110010011110000000001000000000100001000010000000100000000100000000000000000000000000000000000000000000000000000000000000000010001001001001010000000000001011111111000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010010100101010000000000010000000011010110000000010000100001000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000100000001000001000000000000000010110111001000000100000000101010010000100100000001000000000000000000000000000000000000000000000000000000000000000010010001000010000000010000000100000010101101000000000000000010000000000000000001001000010000000000000000000000000000000000000000000000000000001000000000010100010010100001100001010000100110100101000001010000010000001000100001000000000000000000000000000000000000000000000000000000000000000000000000000001000101010100000001101001011110111011010001000000000010000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000010000000010010100001110100000010100100010100000000000010000100001000100100000100000010000000000000000000000000000000000000000000000000000000000000001000000000000000010000110000000000110010001001001010000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000100001010000000101000111011000010000000000010100000010100010001000100000100000010000100000000000000000000000000000000000000000000000000000000000000000000000010000100000000101000000000000000000010000010000000001000010001000000010000100000000000000000000000000000000000000000000100000000000000000000010010000101000010010001000110000000000000000001010001010001001001001001000010000000000000000000000000000000000000000000000010000000000000000000000000010000001010000000001010000010000000000101001001100000000000000100000000000000000000000000000000010000000000000000000000000000000100000000000000000100000110000000100001101000101000000000000000000000010010001010000001010010010100000000000000000000000000000000000000000000000000000000000000000000000010010001000010000100010110011100000000000000000100010000100001001010001000000001001000000000000001000000000000000000000000000000000010000000000000000001000010000001010010101101101000000000000000000000001010010000000010100100000000000000000000001000010000000000100000000000000000100000000001000000000000010101000000000011000000111000000000010000000101010000100101000000100010001000000000010001000010000001000100001000000010000010001010000000000000000000100000100010010100101011010000000000100001000000000010000001000000101001000100000100000000000000000000000000001000000000000001000000000010000100010000010100010000000100101010100000000100101000101100010101010000000001000001000000010001000010100010010000010000000000000010000000100010000001000000000000010000100101010101011010000000000010000010010100010101010010010000101000000000001000010000000010000000000100000010000000010000000001000001000000000000001010000001000001001100000000000001010111011010001000010101000000001010010000000000000001010000100000000000000000100000000101010100000101000000000000000000000000100100110010000000000010001000100000100001010001010001000010000100000101010001000100010000010100000000000000000000000010100000000000000000000000100000010010010000000000000001000101010010011010001010000010101010101001001000001010101010000000000000000001000000000010010000000100000000101010000010000101001010100000000000000000001000000001001001010111010000011010000101001001010010101000000000000000000000000100000001000010010010000000000001000000000001010100000001000000000000000000000000010101100000010101001011100000100110010101101010000000000000000001000001010100100001001001000010100000000000000100000101000000000000000000000000000000010101010010000000101010110100001001010100101000000000010101000000001000000010100001000101010000001000010000010010100000000000101000000000000000000000001000101001000010101111101001010101110101000010000000000000000000100000000000010100101001110000000000000100100100001010000000000000000000000000000000001100100100100000001111101010100101010101010001000000000101001000000101000000100000010101011100000100000100101010101010000000001000000000000000000000000110110101000010010101111010000011111000000000000000001000000010100000010001001001001101111111100001001001010100010101000000000000000000000000000010000010010000001000001010111011101000001101000000000000000000010000001010001001001010101111011111111000100101001000010101100000000100000000000000000000000010101010100000000011111010000000110010010001000001101001000000000000100010001000110111111011111110001001000001011110000000000000000000000000000000000011010100100101001001011111110100001010000100100000000000010001001000000101000101011001011111111111101100000000010111100000000000000000000000000000000000101001001000000101110110100001000100001000010101000010001000000000100000101001101111101111011011110001001000111010100000000000000000000000000000000001001110100010000010011111101000101000000100000001001001000101010010000100001001011111111111111111111000000010001111110000000000000000000000000000000000010101010000000001011111010010000010001000010000100000000000000001010000101010110111111111111111100000000000111010110000000000000000000000000000000000011111010100001010011111111110101000001010000000101001001010000100001010010110110111110111111111111000000001001101111000000000000000000000000000001000000010101000010101011111110010000010100001000101001010010001000000100010010010111111111111111111111000000100111111010000000000000000000000000000000000000011001010100110010101011000001000101000000000000000100001010000001010010001011011111111111111110100000001010101111000000000000000000000000000000000000000010001010011111111100101010010000000100100001000001000001010100001010100111111111111111101111000001011111111011000000000000000000000000001000000000000000000101011011010110101000010000000000001000000000100001000101001010110001111011111111111111011100101111011011000000000000000000000000100010000000000000000100111101011010100001001000100000000000001010011001010001010010000101111111110111111111100001011111111101000000000000000000000000110100100100000000000111011110101010010000001000000010000000010010000100001010010010100010111011111011110111111000101111011111000000000000000000000000100101000000000000000010101011111000101010000010100000000001000100001001010000101001011111011111111111111101100000011111110110001000000000000000000000100101100000000000000000001111010100001000010000100000001000100010000000001001001010000011111111111111111111101001001011111111000000000000000000000000010000000000000000000000000111110100100010100001000010101000000100001000000101010000101001111111111111111010110000011111011100000100000000000000000000000000000000000000000000001111010010001000001000100000001001000010000101010000101010010101111111011010111111111100011111111111000000000000000100000000000000000000000000000000000101010100000001010100000100010010100001000000010010001001001111111111111111110110111001011111111110000001000000000000000000000000010000000000000000000000000010100000000000000101001000100000100001000010101000010101011111011111111111010000001101111110000000000000000000000000000000000000000000000000000000001000010001000010100100100001001010001000100010000101001111111010111101111110111000000111101100000000010001000100000000000000101000000000000000000000010010101000000000010000100100100000000010011000100100101011011111101101011110101000000101111100100000000000000010000000000000010000000000000000000000101000010010010000010100010000000000010000000100100010100111111011111011110111110000000011111000000000000000000000000000000001101010000000000000000000010001010001001010000010001000001001000000100010010000101011111111111100111111011010000101111000000000000000000000000000000001000001010000000000000000010100000000010100000000000000000000010100000000010010010110111110111000011111111000000000110000000000000000000000000000000000100100010000100000000000010101000000010101010100000000001000000010101001000010001010110111111111110110101000000000000000000000000000000000000000000000000001010010010000000000000101010010100010100001000010000100100000000000010001000101011111111111101010110000000000100000000000000000000000000011000000000000000000000000000000000010111010101101010000100010000000000000101000010001001000101001111110111010010100000000001000000000000000000000000001000000000000000000010000000000000010000101010101010100010001000000010010000001000100000010010110111011010101000000000000000000000000000000000000000011100000000000000000010000000000000000111101010110100010000000100010000000101000100001000000100010101101010000010000000000000010000000000000000000000000000100000001000000000000000000000001010011010010010100101010001000001001000010000100010001000000011010000010001010000000000100000000000000000000000010000010000000000000000000000000000000001101011010010010000010010001000100001000000001000000101000000000100000000000000000000000000000000000000000000000001010000000000000000000000000000000000101100101001000001010100100010000000000100100001010000001000010000101000000000000000000000000000000000000000000000000000000000000000100000000000000000100101000000100100001010010001001010100100001000001001000100001010100101010000010000010000000000000000000000000000000000000000000000000000000000000000000000001000010010100010100000101010010001010101000100001000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000101001000010010010101001010101010101011010001000000000000100101000100000000000000000000000000000000000000000000000000000000000000000000000000000011010000010101001000101010001010101001010100001010000100010010000000001000001010000000000000000000000000000000000000000000000000000000000000000000000001101101101010101010010010100100101010100110010000100000010001010010100101001000001000000000000000000000000000000000000000000000000000000000000000000000010100010101010010001010101011010101011001001010010101000100001000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000001011010101010010100101001010101001101010000000000101000100101000010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010010101011010101011111101111110110001010100100010100001001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010101101101011001100001111010110110101011001010000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000101010000000000000000010101011010100100001101000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010111011101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100010000000000001000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

	

	begin

	c_clk_divider: process(in_clk_50mhz) 
	begin
		if rising_edge(in_clk_50mhz) then
			clk_divider <= std_logic_vector(unsigned(clk_divider) + 1);
		end if;
	end process;
	
	e_vgaController: VgaController 
	generic map
	(
		pixelFreq => 25_000_000,

		hSync_visibleArea	=> 640,
		hSync_frontPorch => 16,
		hSync_syncPulse => 96,
		hSync_backPorch => 48,

		vSync_visibleArea	=> 480,
		vSync_frontPorch => 10,
		vSync_syncPulse => 2,
		vSync_backPorch => 33	
	)
	port map
	(
		in_clk => clk_divider(0),
		
		out_vgaRGB 	 => out_vgaRGB,
		out_vgaHSync => out_vgaHSync,
		out_vgaVSync => out_vgaVSync,

		out_isDisplaying	=> isDisplaying,
		out_hPos				=> hPos,
		out_vPos				=> vPos,
		in_vgaRGB			=> rgb
	);
	
	process(clk_divider)
	begin
		if rising_edge(clk_divider(0)) and isDisplaying = '1' then
		
			if vPos < 150 and hPos < 150 then
				position <= vPos*150+hPos;
				rgb <= (imgR(position),imgG(position),imgB(position));

			elsif vPos < 150  and hPos >= 150 and hPos < 300 then
				position <= vPos*150+(hPos-150);
				rgb <= (imgR(position),imgR(position),imgR(position));
				
			elsif vPos < 150  and hPos >= 300 and hPos < 450 then
				position <= vPos*150+(hPos-300);
				rgb <= (imgG(position),imgG(position),imgG(position));
				
			elsif vPos < 150  and hPos >= 450 and hPos < 600 then
				position <= vPos*150+(hPos-450);
				rgb <= (imgB(position),imgB(position),imgB(position));
				
			else
				rgb <= "000";
			end if;
		end if;
	end process;

end behaviour;

